//module lfsr(clk, reset, lfsr);
module lfsr_tb();

reg sim_clk, reset;
wire [4:0] lfsr;

lfsr dut (
.clk(sim_clk),
.reset(reset),
.lfsr(lfsr)
);

// simulation for the clk 
 initial begin
    sim_clk = 0; 
    #5
    forever begin
      sim_clk = 1; 
      #5
      sim_clk = 0; 
      #5  
      sim_clk= 0; 
    end
  end

  initial begin
    reset=0;
    #350


  $stop;
end

endmodule 